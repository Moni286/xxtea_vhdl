--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:58:09 02/11/2018
-- Design Name:   
-- Module Name:   C:/Users/HP/Desktop/University/Academics/Capstone/XXTEA/XXTEA/mx_tb.vhd
-- Project Name:  XXTEA
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mx_add
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY mx_tb IS
END mx_tb;
 
ARCHITECTURE behavior OF mx_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mx_add
    PORT(
         z : IN  std_logic_vector(31 downto 0);
         y : IN  std_logic_vector(31 downto 0);
         addend : IN  std_logic_vector(31 downto 0);
         sum : IN  std_logic_vector(31 downto 0);
         key : IN  std_logic_vector(31 downto 0);
         sigma : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal z : std_logic_vector(31 downto 0) := (others => '0');
   signal y : std_logic_vector(31 downto 0) := (others => '0');
   signal addend : std_logic_vector(31 downto 0) := (others => '0');
   signal sum : std_logic_vector(31 downto 0) := (others => '0');
   signal key : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal sigma : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: mx_add PORT MAP (
          z => z,
          y => y,
          addend => addend,
          sum => sum,
          key => key,
          sigma => sigma
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      z <= x"bbbbbbbb";
		y <= x"aaaaaaac";
		addend <= x"cccccccc";
		key <= x"eeeeeeee";
		sum <= x"9e3779b9";
      

      wait;
   end process;

END;
